module main

import strings

// resolve_type_alias resolves type alias chains to the underlying type.
// V doesn't allow type A = B where B is also a type alias.
fn (mut c C2V) resolve_type_alias(type_name string) string {
	// If this type is a known alias, resolve to its underlying type
	if underlying := c.type_aliases[type_name] {
		// Recursively resolve in case of chains
		return c.resolve_type_alias(underlying)
	}
	return type_name
}

// |-RecordDecl 0x7fd7c302c560 <a.c:3:1, line:5:1> line:3:8 struct User definition
fn (mut c C2V) record_decl(node &Node) {
	vprintln('record_decl("${node.name}")')
	// Skip empty structs (extern or forward decls)
	if node.kindof(.record_decl) && node.inner.len == 0 {
		return
	}
	mut c_name := node.name
	// Dont generate struct header if it was already generated by typedef
	// Confusing, but typedefs in C AST are really messy.
	// ...
	// If the struct has no name, then it's `typedef struct { ... } name`
	// AST: 1) RecordDecl struct definition 2) TypedefDecl struct name
	if c.tree.inner.len > c.node_i + 1 {
		next_node := c.tree.inner[c.node_i + 1]
		if next_node.kind == .typedef_decl {
			if c.is_verbose {
				c.genln('// typedef struct')
			}
			c_name = next_node.name
			if c_name.contains('apthing_t') {
				vprintln(node.str())
			}
		}
	}

	if c_name in builtin_type_names {
		return
	}
	if c.is_verbose {
		c.genln('// struct decl name="${c_name}"')
	}
	if c_name in c.types {
		if node.previous_declaration == '' {
			return
		}
	}
	// Anonymous struct, most likely the next node is a vardecl with this anon struct type, so remember it
	if c_name == '' {
		c_name = 'AnonStruct_${node.location.line}'
		c.last_declared_type_name = c_name
	}

	// First pass: scan for anonymous enums and generate named enum types BEFORE the struct.
	// V doesn't support inline `enum {}` in struct fields like it does for struct/union.
	// We need to generate the enum as a separate named type.
	mut anon_enum_names := map[int]string{} // maps field index to generated enum name
	mut struct_v_name := c.add_struct_name(mut c.types, c_name)
	mut pending_enum := &Node(unsafe { nil })
	for i, field in node.inner {
		if field.kind == .enum_decl {
			pending_enum = unsafe { &node.inner[i] }
			continue
		}
		if field.kind == .field_decl && pending_enum != unsafe { nil } {
			field_type := convert_type(field.ast_type.qualified)
			if field_type.name.contains('unnamed enum at') {
				// Generate a named enum for this anonymous enum
				field_name := filter_name(field.name, false)
				enum_name := c.generate_named_enum_for_anon(pending_enum, struct_v_name, field_name)
				anon_enum_names[i] = enum_name
			}
			pending_enum = unsafe { nil }
		}
	}

	if c_name !in ['struct', 'union'] {
		// prevent duplicate generations:
		if struct_v_name in c.generated_declarations {
			return
		}
		c.generated_declarations[struct_v_name] = true
		if node.tags.contains('union') {
			c.genln('union ${struct_v_name} { ')
		} else {
			c.genln('struct ${struct_v_name} { ')
		}
	}
	mut new_struct := Struct{}
	// in V it's `field struct {...}`, but in C we get struct definition first, so save it and use it in the
	// next child
	mut anon_struct_definition := ''
	mut anon_enum_definition := ''
	for i, field in node.inner {
		c.gen_comment(field)
		// Handle anon structs and unions (unions appear as RecordDecl with tagUsed='union')
		if field.kind == .record_decl {
			is_union := field.tags.contains('union')
			anon_struct_definition = c.anon_struct_field_type(field, is_union)
			continue
		}
		if field.kind == .union_decl {
			anon_struct_definition = c.anon_struct_field_type(field, true)
			continue
		}
		// Handle anon enums - skip, already processed in first pass
		if field.kind == .enum_decl {
			continue
		}
		// There may be comments, skip them
		if field.kind != .field_decl {
			continue
		}
		field_type := convert_type(field.ast_type.qualified)
		filtered := filter_name(field.name, false)
		// Don't uncapitalize if it's a C. prefixed name (builtin function)
		field_name := if filtered.starts_with('C.') { filtered[2..] + '_' } else { filtered.uncapitalize() }
		mut field_type_name := field_type.name

		// Handle anon structs/unions, the anonymous type has just been defined above, use its definition
		// Note: "unnamed struct at" and "unnamed union at" both need to be handled
		if (field_type_name.contains('unnamed struct at') || field_type_name.contains('unnamed union at') || field_type_name.contains('(unnamed at')) && !field_type_name.contains('unnamed enum') {
			field_type_name = anon_struct_definition
		}
		// Handle anon enums - use the pre-generated named enum type
		if field_type_name.contains('unnamed enum at') {
			if i in anon_enum_names {
				field_type_name = anon_enum_names[i]
			} else {
				field_type_name = anon_enum_definition
			}
		}
		if field_type_name.contains('anonymous at') {
			continue
		}
		/*
		if field_type.name.contains('union') {
			continue // TODO
		}
		*/
		new_struct.fields << field_name
		if field_type.name.ends_with('_s') { // TODO doom _t _s hack, remove
			n := field_type.name[..field_type.name.len - 2] + '_t'
			c.genln('\t${field_name} ${c.prefix_external_type(n)}')
		} else {
			c.genln('\t${field_name} ${c.prefix_external_type(field_type_name)}')
		}
	}
	c.structs[c_name] = new_struct
	c.genln('}')
}

fn (mut c C2V) anon_struct_field_type(node &Node, is_union bool) string {
	mut sb := strings.new_builder(50)
	if is_union {
		sb.write_string('union {\n')
	} else {
		sb.write_string('struct {\n')
	}
	mut nested_anon_def := ''
	for field in node.inner {
		// Handle nested anonymous struct/union definitions
		if field.kind == .record_decl {
			nested_is_union := field.tags.contains('union')
			nested_anon_def = c.anon_struct_field_type(field, nested_is_union)
			continue
		}
		if field.kind != .field_decl {
			continue
		}
		field_type := convert_type(field.ast_type.qualified)
		field_name := filter_name(field.name, false)
		mut field_type_name := field_type.name
		// Use nested anonymous definition if this field references one
		if field_type_name.contains('unnamed struct at') || field_type_name.contains('unnamed union at') || field_type_name.contains('(unnamed at') || field_type_name.contains('anonymous at') {
			field_type_name = nested_anon_def
		}
		// Apply external type prefix for types from headers
		field_type_name = c.prefix_external_type(field_type_name)
		sb.write_string('${field_name} ${field_type_name}\n')
	}
	sb.write_string('}')
	return sb.str()
}

fn (mut c C2V) anon_enum_field_type(node &Node) string {
	mut sb := strings.new_builder(50)
	sb.write_string('enum {\n')
	for i, child in node.inner {
		if child.kind != .enum_constant_decl {
			continue
		}
		c_name := filter_name(child.name, false)
		v_name := c_name.camel_to_snake().trim_left('_')
		sb.write_string('${v_name}')
		// handle custom enum vals, e.g. `MF_SHOOTABLE = 4`
		if child.inner.len > 0 {
			mut const_expr := child.inner[0]
			if const_expr.kind == .constant_expr && const_expr.inner.len > 0 {
				// Try to get the literal value
				literal := const_expr.inner[0]
				if literal.kind == .integer_literal {
					sb.write_string(' = ${literal.value.to_str()}')
				}
			}
		}
		sb.write_string('\n')
		_ = i
	}
	sb.write_string('}')
	return sb.str()
}

// Generate a named enum type for an anonymous enum field in a struct.
// V doesn't support inline `enum {}` syntax in struct fields (unlike struct/union),
// so we generate a separate named enum type before the struct.
// Returns the generated enum type name.
fn (mut c C2V) generate_named_enum_for_anon(node &Node, struct_name string, field_name string) string {
	// Create enum name from struct name + field name, e.g. "With_anon_enum_Status"
	enum_name := '${struct_name}_${field_name.capitalize()}'

	// Generate the enum definition
	c.genln('enum ${enum_name} {')
	for child in node.inner {
		if child.kind != .enum_constant_decl {
			continue
		}
		c_name := filter_name(child.name, false)
		v_name := c_name.camel_to_snake().trim_left('_')
		mut line := '\t${v_name}'
		// handle custom enum vals, e.g. `MF_SHOOTABLE = 4`
		if child.inner.len > 0 {
			mut const_expr := child.inner[0]
			if const_expr.kind == .constant_expr && const_expr.inner.len > 0 {
				// Try to get the literal value
				literal := const_expr.inner[0]
				if literal.kind == .integer_literal {
					line += ' = ${literal.value.to_str()}'
				}
			}
		}
		c.genln(line)
	}
	c.genln('}')
	c.genln('')

	return enum_name
}

// Typedef node goes after struct enum, but we need to parse it first, so that "type name { " is
// generated first
fn (mut c C2V) typedef_decl(node &Node) {
	mut typ := node.ast_type.qualified
	// just a single line typedef: (alias)
	// typedef sha1_context_t sha1_context_s ;
	// typedef after enum decl, just generate "enum NAME {" header
	mut c_alias_name := node.name // get_val(-2)
	if c_alias_name.contains('et_context_t') {
		// TODO remove this
		return
	}
	if c_alias_name in builtin_type_names {
		return
	}

	if c_alias_name in c.types || c_alias_name in c.enums {
		// This means that this is a struct/enum typedef that has already been defined.
		return
	}

	v_alias_name := c.add_struct_name(mut c.types, c_alias_name)

	if typ.starts_with('struct ') && typ.ends_with(' *') {
		// Opaque pointer, for example: typedef struct TSTexture_t *TSTexture;
		c.genln('type ${v_alias_name} = voidptr')
		return
	}

	if !typ.contains(c_alias_name) {
		// Function pointer: int (*)(args)
		if typ.contains('(*)') {
			tt := convert_type(typ)
			typ = c.prefix_external_type(tt.name)
		}
		// Function type without pointer: int (args) - e.g., typedef int fn_name(args)
		// Note: don't require comma - single-argument functions like "void (void *)" have no comma
		else if typ.contains('(') && typ.contains(')') && !typ.starts_with('(') {
			// Parse function type: "int (arg1, arg2, ...)" -> "fn (arg1, arg2) int"
			ret_typ := convert_type(typ.all_before('(').trim_space())
			mut s := 'fn ('
			sargs := typ.find_between('(', ')')
			args := sargs.split(',')
			for i, arg in args {
				t := convert_type(arg.trim_space())
				s += c.prefix_external_type(t.name)
				if i < args.len - 1 {
					s += ', '
				}
			}
			if ret_typ.name == 'void' {
				typ = s + ')'
			} else {
				typ = '${s}) ${c.prefix_external_type(ret_typ.name)}'
			}
			typ = typ.replace('(void)', '()')
		}
		// Struct types have junk before spaces
		else {
			c_alias_name = c_alias_name.all_after(' ')
			tt := convert_type(typ)
			typ = c.prefix_external_type(tt.name)
		}
		if c_alias_name.starts_with('__') {
			// Skip internal stuff like __builtin_ms_va_list
			return
		}
		if typ in c.enums {
			return
		}

		mut cgen_alias := typ
		if cgen_alias.starts_with('_') {
			cgen_alias = trim_underscores(typ)
		}
		if typ !in ['int', 'i8', 'i16', 'i64', 'u8', 'u16', 'u32', 'u64', 'f32', 'f64', 'usize', 'isize', 'bool', 'void', 'voidptr']
			&& !typ.starts_with('fn (') {
			// TODO handle this better
			cgen_alias = cgen_alias.capitalize()
		}
		// Resolve type alias chains - V doesn't allow type A = B where B is an alias
		resolved_alias := c.resolve_type_alias(cgen_alias)
		prefixed_alias := c.prefix_external_type(resolved_alias)
		// Store this alias mapping for future resolution
		c.type_aliases[c_alias_name.capitalize()] = prefixed_alias
		c.genln('type ${c_alias_name.capitalize()} = ${prefixed_alias}') // typedef alias (SINGLE LINE)')
		return
	}
	if typ.contains('enum ') {
		// enums were alredy handled in enum_decl
		return
	} else if typ.contains('struct ') {
		// structs were already handled in struct_decl
		return
	} else if typ.contains('union ') {
		// unions were alredy handled in struct_decl
		return
	}
}

// this calls typedef_decl() above
fn (mut c C2V) parse_next_typedef() bool {
	// Hack: typedef with the actual enum name is next, parse it and generate "enum NAME {" first
	/*
	XTODO
	next_line := c.lines[c.line_i + 1]
	if next_line.contains('TypedefDecl') {
		c.line_i++
		c.parse_next_node()
		return true
	}
	*/
	return false
}
